module L2part6(s,u,v,w,x,y,m0,m1,m2,m3,m4,m5,m6,m7 ,led,HEX0, HEX1, HEX2, HEX3, HEX4,HEX5,HEX6,HEX7);

	input [2:0]s,u,v,w,x,y;
	
   output [0:6]HEX0, HEX1, HEX2, HEX3, HEX4, HEX5, HEX6, HEX7;
   output [2:0]m0,m1,m2,m3,m4,m5,m6,m7;
   output [17:0]led;
   
   assign led[17:15] = s;
	assign led[14:12] = u;
	assign led[11:9] = v;
	assign led[8:6] = w;
	assign led[5:3] = x;
	assign led[2:0] = y;
   
	assign m7 =  (s ==3'b011) ? u :
               (s ==3'b100) ? v :
               (s ==3'b101) ? w :
               (s ==3'b110) ? w :
					(s ==3'b111) ? x :y;
					
	assign m6 =  (s ==3'b010) ? u :
               (s ==3'b011) ? v :
               (s ==3'b100) ? w :
               (s ==3'b101) ? w :
					(s ==3'b110) ? x :y;
					
	assign m5 =  (s ==3'b001) ? u :
               (s ==3'b010) ? v :
               (s ==3'b011) ? w :
               (s ==3'b100) ? w :
					(s ==3'b101) ? x :y;	
								
   assign m4 =  (s ==3'b000) ? u :
               (s ==3'b001) ? v :
               (s ==3'b010) ? w :
               (s ==3'b011) ? w :
					(s ==3'b100) ? x :y;
               
   assign m3 =  (s ==3'b000) ? v :
               (s ==3'b001) ? w :
               (s ==3'b010) ? w :
               (s ==3'b011) ? x :
					(s ==3'b111) ? u : y;
               
   assign m2 =  (s ==3'b000) ? w :
               (s ==3'b001) ? w :
               (s ==3'b010) ? x :
               (s ==3'b110) ? u :
					(s ==3'b111) ? v : y;
               
   assign m1 =  (s ==3'b000) ? w :
               (s ==3'b001) ? x :
               (s ==3'b101) ? u :
               (s ==3'b110) ? v :
					(s ==3'b111) ? w : y;
				
               
   assign m0 =  (s ==3'b000) ? x :
               (s ==3'b100) ? u :
               (s ==3'b101) ? v :
               (s ==3'b110) ? w :
					(s ==3'b111) ? w : y;
               
	assign HEX7 = (m7 ==3'b000) ? 7'b1001000:
                 (m7 ==3'b001) ? 7'b0110000:
                 (m7 ==3'b010) ? 7'b1110001:
                 (m7 ==3'b011) ? 7'b0000001: 7'b1111111;
					  
	assign HEX6 = (m6 ==3'b000) ? 7'b1001000:
                 (m6 ==3'b001) ? 7'b0110000:
                 (m6 ==3'b010) ? 7'b1110001:
                 (m6 ==3'b011) ? 7'b0000001: 7'b1111111;
					  
	assign HEX5 = (m5 ==3'b000) ? 7'b1001000:
                 (m5 ==3'b001) ? 7'b0110000:
                 (m5 ==3'b010) ? 7'b1110001:
                 (m5 ==3'b011) ? 7'b0000001: 7'b1111111;
   
   assign HEX4 = (m4 ==3'b000) ? 7'b1001000:
                 (m4 ==3'b001) ? 7'b0110000:
                 (m4 ==3'b010) ? 7'b1110001:
                 (m4 ==3'b011) ? 7'b0000001: 7'b1111111;
                 
   assign HEX3 = (m3 ==3'b000) ? 7'b1001000:
                 (m3 ==3'b001) ? 7'b0110000:
                 (m3 ==3'b010) ? 7'b1110001:
                 (m3 ==3'b011) ? 7'b0000001: 7'b1111111;
                 
   assign HEX2 = (m2 ==3'b000) ? 7'b1001000:
                 (m2 ==3'b001) ? 7'b0110000:
                 (m2 ==3'b010) ? 7'b1110001:
                 (m2 ==3'b011) ? 7'b0000001: 7'b1111111;
                 
                 
   assign HEX1 = (m1 ==3'b000) ? 7'b1001000:
                 (m1 ==3'b001) ? 7'b0110000:
                 (m1 ==3'b010) ? 7'b1110001:
                 (m1 ==3'b011) ? 7'b0000001: 7'b1111111;
                 
   assign HEX0 = (m0 ==3'b000) ? 7'b1001000:
                 (m0 ==3'b001) ? 7'b0110000:
                 (m0 ==3'b010) ? 7'b1110001:
                 (m0 ==3'b011) ? 7'b0000001: 7'b1111111;

endmodule
