module ledtest(sw,ledr);

	input [2:0]sw;
	output [2:0]ledr;
	
	assign ledr=sw;
	
endmodule
