module not_gate(A1,out);

input A1;
output out;
assign out=~A1;

endmodule
